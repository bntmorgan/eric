`define CSR_DDR3_CSR_CTRL 10'h000
`define CSR_DDR3_CSR_STAT 10'h001
`define CSR_DDR3_CSR_ADDR 10'h002
`define CSR_DDR3_CSR_W0 10'h003
`define CSR_DDR3_CSR_W1 10'h004
`define CSR_DDR3_CSR_W2 10'h005
`define CSR_DDR3_CSR_W3 10'h006
`define CSR_DDR3_CSR_W4 10'h007
`define CSR_DDR3_CSR_W5 10'h008
`define CSR_DDR3_CSR_W6 10'h009
`define CSR_DDR3_CSR_W7 10'h00a
`define CSR_DDR3_CSR_R0 10'h00b
`define CSR_DDR3_CSR_R1 10'h00c
`define CSR_DDR3_CSR_R2 10'h00d
`define CSR_DDR3_CSR_R3 10'h00e
`define CSR_DDR3_CSR_R4 10'h00f
`define CSR_DDR3_CSR_R5 10'h010
`define CSR_DDR3_CSR_R6 10'h011
`define CSR_DDR3_CSR_R7 10'h012
`define CSR_DDR3_CSR_GWTC 10'h013
`define CSR_DDR3_CSR_GRTC 10'h014
