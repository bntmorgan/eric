`ifndef __TRN_VH__
`define __TRN_VH__

`define TRN_CSR_STAT_TRN          10'h000
`define TRN_CSR_CFG_PCI_ADDR      10'h001
`define TRN_CSR_CFG_COMMAND       10'h002
`define TRN_CSR_CFG_DSTATUS       10'h003
`define TRN_CSR_CFG_DCOMMAND      10'h004
`define TRN_CSR_CFG_DCOMMAND2     10'h005
`define TRN_CSR_CFG_LSTATUS       10'h006
`define TRN_CSR_CFG_LCOMMAND      10'h007
`define TRN_CSR_TRN_FC_CPLD       10'h008
`define TRN_CSR_TRN_FC_CPLH       10'h009
`define TRN_CSR_TRN_FC_NPD        10'h00a
`define TRN_CSR_TRN_FC_NPH        10'h00b
`define TRN_CSR_TRN_FC_PD         10'h00c
`define TRN_CSR_TRN_FC_PH         10'h00d
`define TRN_CSR_TRN_FC_SEL        10'h00e

`endif//__TRN_VH__
