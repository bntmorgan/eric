module mpu_decoder (
  // Instruction to decode
);

endmodule
