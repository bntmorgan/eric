/**
 * 30.000% Makina Process Unit
 */

`define MPU_OP_MASK   4'h1
`define MPU_OP_CMP    4'h2
`define MPU_OP_LT     4'h3
`define MPU_OP_ADD    4'h4
`define MPU_OP_INT    4'hc
`define MPU_OP_MLOAD  4'hd
`define MPU_OP_LOAD   4'he
`define MPU_OP_JMP    4'hf
