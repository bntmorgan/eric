module main();

initial begin
  $finish();
end

endmodule
